/*
Author: Ganesg
Date : 01/12/2024

*/

//Instruction Memory

module Instruction_Mem(
	input clk,
	input reset,
	input [31:0] read_address,
	output [31:0] instruction_out
);

re


endmodule