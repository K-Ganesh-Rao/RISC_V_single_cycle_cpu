/*
Author: Ganesg
Date : 01/12/2024

*/

//Register file

module Reg_file